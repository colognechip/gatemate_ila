library ieee;
use ieee.std_logic_1164.all;

package const_image is
 constant CLKFRQ           : integer := 10_000_000;
 end const_image;
